module memoryBank (mem_data_out,mem_data_in,mem_addr_out,mem_addr_in,enable,reset);
output reg [7:0] mem_data_out;
input [7:0] mem_data_in;
input [4:0] mem_addr_in,mem_addr_out;
input enable,reset;



endmodule //memoryBank